/******************************************************************************

    File Name:  COREPWM.v
      Version:  4.0
         Date:  July 20th, 2009
  Description:  Top level module
  
  
  SVN Revision Information:
  SVN $Revision: 10267 $
  SVN $Date: 2009-10-15 16:42:37 -0700 (Thu, 15 Oct 2009) $  
  
  

 COPYRIGHT 2009 BY ACTEL 
 THE INFORMATION CONTAINED IN THIS DOCUMENT IS SUBJECT TO LICENSING RESTRICTIONS 
 FROM ACTEL CORP.  IF YOU ARE NOT IN POSSESSION OF WRITTEN AUTHORIZATION FROM 
 ACTEL FOR USE OF THIS FILE, THEN THE FILE SHOULD BE IMMEDIATELY DESTROYED AND 
 NO BACK-UP OF THE FILE SHOULD BE MADE. 
 
FUNCTIONAL DESCRIPTION:  
Refer to the CorePWM Handbook.
******************************************************************************/
`timescale 1ns/1ns
module
corepwm
#
(
parameter
FAMILY
=
0
,
parameter
CONFIG_MODE
=
0
,
parameter
PWM_NUM
=
1
,
parameter
APB_DWIDTH
=
8
,
parameter
FIXED_PRESCALE_EN
=
1
,
parameter
FIXED_PRESCALE
=
8
,
parameter
FIXED_PERIOD_EN
=
0
,
parameter
FIXED_PERIOD
=
8
,
parameter
DAC_MODE1
=
0
,
parameter
DAC_MODE2
=
0
,
parameter
DAC_MODE3
=
0
,
parameter
DAC_MODE4
=
0
,
parameter
DAC_MODE5
=
0
,
parameter
DAC_MODE6
=
0
,
parameter
DAC_MODE7
=
0
,
parameter
DAC_MODE8
=
0
,
parameter
DAC_MODE9
=
0
,
parameter
DAC_MODE10
=
0
,
parameter
DAC_MODE11
=
0
,
parameter
DAC_MODE12
=
0
,
parameter
DAC_MODE13
=
0
,
parameter
DAC_MODE14
=
0
,
parameter
DAC_MODE15
=
0
,
parameter
DAC_MODE16
=
0
,
parameter
SHADOW_REG_EN1
=
0
,
parameter
SHADOW_REG_EN2
=
0
,
parameter
SHADOW_REG_EN3
=
0
,
parameter
SHADOW_REG_EN4
=
0
,
parameter
SHADOW_REG_EN5
=
0
,
parameter
SHADOW_REG_EN6
=
0
,
parameter
SHADOW_REG_EN7
=
0
,
parameter
SHADOW_REG_EN8
=
0
,
parameter
SHADOW_REG_EN9
=
0
,
parameter
SHADOW_REG_EN10
=
0
,
parameter
SHADOW_REG_EN11
=
0
,
parameter
SHADOW_REG_EN12
=
0
,
parameter
SHADOW_REG_EN13
=
0
,
parameter
SHADOW_REG_EN14
=
0
,
parameter
SHADOW_REG_EN15
=
0
,
parameter
SHADOW_REG_EN16
=
0
,
parameter
FIXED_PWM_POS_EN1
=
1
,
parameter
FIXED_PWM_POS_EN2
=
1
,
parameter
FIXED_PWM_POS_EN3
=
1
,
parameter
FIXED_PWM_POS_EN4
=
1
,
parameter
FIXED_PWM_POS_EN5
=
1
,
parameter
FIXED_PWM_POS_EN6
=
1
,
parameter
FIXED_PWM_POS_EN7
=
1
,
parameter
FIXED_PWM_POS_EN8
=
1
,
parameter
FIXED_PWM_POS_EN9
=
1
,
parameter
FIXED_PWM_POS_EN10
=
1
,
parameter
FIXED_PWM_POS_EN11
=
1
,
parameter
FIXED_PWM_POS_EN12
=
1
,
parameter
FIXED_PWM_POS_EN13
=
1
,
parameter
FIXED_PWM_POS_EN14
=
1
,
parameter
FIXED_PWM_POS_EN15
=
1
,
parameter
FIXED_PWM_POS_EN16
=
1
,
parameter
FIXED_PWM_POSEDGE1
=
0
,
parameter
FIXED_PWM_POSEDGE2
=
0
,
parameter
FIXED_PWM_POSEDGE3
=
0
,
parameter
FIXED_PWM_POSEDGE4
=
0
,
parameter
FIXED_PWM_POSEDGE5
=
0
,
parameter
FIXED_PWM_POSEDGE6
=
0
,
parameter
FIXED_PWM_POSEDGE7
=
0
,
parameter
FIXED_PWM_POSEDGE8
=
0
,
parameter
FIXED_PWM_POSEDGE9
=
0
,
parameter
FIXED_PWM_POSEDGE10
=
0
,
parameter
FIXED_PWM_POSEDGE11
=
0
,
parameter
FIXED_PWM_POSEDGE12
=
0
,
parameter
FIXED_PWM_POSEDGE13
=
0
,
parameter
FIXED_PWM_POSEDGE14
=
0
,
parameter
FIXED_PWM_POSEDGE15
=
0
,
parameter
FIXED_PWM_POSEDGE16
=
0
,
parameter
FIXED_PWM_NEG_EN1
=
0
,
parameter
FIXED_PWM_NEG_EN2
=
0
,
parameter
FIXED_PWM_NEG_EN3
=
0
,
parameter
FIXED_PWM_NEG_EN4
=
0
,
parameter
FIXED_PWM_NEG_EN5
=
0
,
parameter
FIXED_PWM_NEG_EN6
=
0
,
parameter
FIXED_PWM_NEG_EN7
=
0
,
parameter
FIXED_PWM_NEG_EN8
=
0
,
parameter
FIXED_PWM_NEG_EN9
=
0
,
parameter
FIXED_PWM_NEG_EN10
=
0
,
parameter
FIXED_PWM_NEG_EN11
=
0
,
parameter
FIXED_PWM_NEG_EN12
=
0
,
parameter
FIXED_PWM_NEG_EN13
=
0
,
parameter
FIXED_PWM_NEG_EN14
=
0
,
parameter
FIXED_PWM_NEG_EN15
=
0
,
parameter
FIXED_PWM_NEG_EN16
=
0
,
parameter
FIXED_PWM_NEGEDGE1
=
0
,
parameter
FIXED_PWM_NEGEDGE2
=
0
,
parameter
FIXED_PWM_NEGEDGE3
=
0
,
parameter
FIXED_PWM_NEGEDGE4
=
0
,
parameter
FIXED_PWM_NEGEDGE5
=
0
,
parameter
FIXED_PWM_NEGEDGE6
=
0
,
parameter
FIXED_PWM_NEGEDGE7
=
0
,
parameter
FIXED_PWM_NEGEDGE8
=
0
,
parameter
FIXED_PWM_NEGEDGE9
=
0
,
parameter
FIXED_PWM_NEGEDGE10
=
0
,
parameter
FIXED_PWM_NEGEDGE11
=
0
,
parameter
FIXED_PWM_NEGEDGE12
=
0
,
parameter
FIXED_PWM_NEGEDGE13
=
0
,
parameter
FIXED_PWM_NEGEDGE14
=
0
,
parameter
FIXED_PWM_NEGEDGE15
=
0
,
parameter
FIXED_PWM_NEGEDGE16
=
0
,
parameter
PWM_STRETCH_VALUE1
=
0
,
parameter
PWM_STRETCH_VALUE2
=
0
,
parameter
PWM_STRETCH_VALUE3
=
0
,
parameter
PWM_STRETCH_VALUE4
=
0
,
parameter
PWM_STRETCH_VALUE5
=
0
,
parameter
PWM_STRETCH_VALUE6
=
0
,
parameter
PWM_STRETCH_VALUE7
=
0
,
parameter
PWM_STRETCH_VALUE8
=
0
,
parameter
PWM_STRETCH_VALUE9
=
0
,
parameter
PWM_STRETCH_VALUE10
=
0
,
parameter
PWM_STRETCH_VALUE11
=
0
,
parameter
PWM_STRETCH_VALUE12
=
0
,
parameter
PWM_STRETCH_VALUE13
=
0
,
parameter
PWM_STRETCH_VALUE14
=
0
,
parameter
PWM_STRETCH_VALUE15
=
0
,
parameter
PWM_STRETCH_VALUE16
=
0
,
parameter
TACH_NUM
=
1
,
parameter
TACH_EDGE1
=
0
,
parameter
TACH_EDGE2
=
0
,
parameter
TACH_EDGE3
=
0
,
parameter
TACH_EDGE4
=
0
,
parameter
TACH_EDGE5
=
0
,
parameter
TACH_EDGE6
=
0
,
parameter
TACH_EDGE7
=
0
,
parameter
TACH_EDGE8
=
0
,
parameter
TACH_EDGE9
=
0
,
parameter
TACH_EDGE10
=
0
,
parameter
TACH_EDGE11
=
0
,
parameter
TACH_EDGE12
=
0
,
parameter
TACH_EDGE13
=
0
,
parameter
TACH_EDGE14
=
0
,
parameter
TACH_EDGE15
=
0
,
parameter
TACH_EDGE16
=
0
,
parameter
TACHINT_ACT_LEVEL
=
0
)
(
input
PRESETN,
input
PCLK,
input
PSEL,
input
PENABLE,
input
PWRITE,
input
[
7
:
0
]
PADDR,
input
[
APB_DWIDTH
-
1
:
0
]
PWDATA,
output
[
APB_DWIDTH
-
1
:
0
]
PRDATA,
output
PREADY,
output
PSLVERR,
input
[
TACH_NUM
-
1
:
0
]
TACHIN,
output
TACHINT,
output
[
PWM_NUM
:
1
]
PWM
)
;
wire
[
APB_DWIDTH
-
1
:
0
]
prescale_reg
,
period_reg
,
period_cnt
;
wire
[
PWM_NUM
:
1
]
pwm_enable_reg
;
wire
[
PWM_NUM
*
APB_DWIDTH
:
1
]
pwm_posedge_reg
,
pwm_negedge_reg
;
wire
sync_pulse
;
wire
[
PWM_NUM
:
1
]
CPWMO
;
reg
[
15
:
0
]
CPWMI
;
wire
[
PWM_NUM
-
1
:
0
]
CPWMl
;
wire
[
TACH_NUM
-
1
:
0
]
TACH_EDGE
;
wire
CPWMOI
;
reg
[
3
:
0
]
CPWMII
;
reg
[
PWM_NUM
-
1
:
0
]
PWM_STRETCH
;
reg
[
TACH_NUM
-
1
:
0
]
CPWMlI
;
reg
[
TACH_NUM
-
1
:
0
]
TACHMODE
;
reg
[
TACH_NUM
-
1
:
0
]
TACHSTATUS
;
reg
[
10
:
0
]
CPWMOl
;
reg
[
10
:
0
]
CPWMIl
;
reg
[
10
:
0
]
CPWMll
;
reg
tach_cnt_clk
;
wire
[
15
:
0
]
TACHPULSEDUR
[
TACH_NUM
-
1
:
0
]
;
wire
[
TACH_NUM
-
1
:
0
]
update_status
;
reg
[
TACH_NUM
-
1
:
0
]
status_clear
;
wire
[
APB_DWIDTH
-
1
:
0
]
CPWMO0
;
parameter
[
15
:
0
]
all_ones
=
16
'h
ffff
;
parameter
[
15
:
0
]
DAC_MODE
=
(
DAC_MODE16
<<
15
)
|
(
DAC_MODE15
<<
14
)
|
(
DAC_MODE14
<<
13
)
|
(
DAC_MODE13
<<
12
)
|
(
DAC_MODE12
<<
11
)
|
(
DAC_MODE11
<<
10
)
|
(
DAC_MODE10
<<
9
)
|
(
DAC_MODE9
<<
8
)
|
(
DAC_MODE8
<<
7
)
|
(
DAC_MODE7
<<
6
)
|
(
DAC_MODE6
<<
5
)
|
(
DAC_MODE5
<<
4
)
|
(
DAC_MODE4
<<
3
)
|
(
DAC_MODE3
<<
2
)
|
(
DAC_MODE2
<<
1
)
|
(
DAC_MODE1
<<
0
)
;
parameter
[
15
:
0
]
SHADOW_REG_EN
=
(
SHADOW_REG_EN16
<<
15
)
|
(
SHADOW_REG_EN15
<<
14
)
|
(
SHADOW_REG_EN14
<<
13
)
|
(
SHADOW_REG_EN13
<<
12
)
|
(
SHADOW_REG_EN12
<<
11
)
|
(
SHADOW_REG_EN11
<<
10
)
|
(
SHADOW_REG_EN10
<<
9
)
|
(
SHADOW_REG_EN9
<<
8
)
|
(
SHADOW_REG_EN8
<<
7
)
|
(
SHADOW_REG_EN7
<<
6
)
|
(
SHADOW_REG_EN6
<<
5
)
|
(
SHADOW_REG_EN5
<<
4
)
|
(
SHADOW_REG_EN4
<<
3
)
|
(
SHADOW_REG_EN3
<<
2
)
|
(
SHADOW_REG_EN2
<<
1
)
|
(
SHADOW_REG_EN1
<<
0
)
;
parameter
[
15
:
0
]
FIXED_PWM_POS_EN
=
(
FIXED_PWM_POS_EN16
<<
15
)
|
(
FIXED_PWM_POS_EN15
<<
14
)
|
(
FIXED_PWM_POS_EN14
<<
13
)
|
(
FIXED_PWM_POS_EN13
<<
12
)
|
(
FIXED_PWM_POS_EN12
<<
11
)
|
(
FIXED_PWM_POS_EN11
<<
10
)
|
(
FIXED_PWM_POS_EN10
<<
9
)
|
(
FIXED_PWM_POS_EN9
<<
8
)
|
(
FIXED_PWM_POS_EN8
<<
7
)
|
(
FIXED_PWM_POS_EN7
<<
6
)
|
(
FIXED_PWM_POS_EN6
<<
5
)
|
(
FIXED_PWM_POS_EN5
<<
4
)
|
(
FIXED_PWM_POS_EN4
<<
3
)
|
(
FIXED_PWM_POS_EN3
<<
2
)
|
(
FIXED_PWM_POS_EN2
<<
1
)
|
(
FIXED_PWM_POS_EN1
<<
0
)
;
parameter
[
15
:
0
]
FIXED_PWM_NEG_EN
=
(
FIXED_PWM_NEG_EN16
<<
15
)
|
(
FIXED_PWM_NEG_EN15
<<
14
)
|
(
FIXED_PWM_NEG_EN14
<<
13
)
|
(
FIXED_PWM_NEG_EN13
<<
12
)
|
(
FIXED_PWM_NEG_EN12
<<
11
)
|
(
FIXED_PWM_NEG_EN11
<<
10
)
|
(
FIXED_PWM_NEG_EN10
<<
9
)
|
(
FIXED_PWM_NEG_EN9
<<
8
)
|
(
FIXED_PWM_NEG_EN8
<<
7
)
|
(
FIXED_PWM_NEG_EN7
<<
6
)
|
(
FIXED_PWM_NEG_EN6
<<
5
)
|
(
FIXED_PWM_NEG_EN5
<<
4
)
|
(
FIXED_PWM_NEG_EN4
<<
3
)
|
(
FIXED_PWM_NEG_EN3
<<
2
)
|
(
FIXED_PWM_NEG_EN2
<<
1
)
|
(
FIXED_PWM_NEG_EN1
<<
0
)
;
parameter
[
16
*
APB_DWIDTH
-
1
:
0
]
FIXED_PWM_POSEDGE
=
{
FIXED_PWM_POSEDGE16
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE15
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE14
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE13
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE12
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE11
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE10
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE9
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE8
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE7
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE6
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE5
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE4
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE3
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE2
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_POSEDGE1
[
APB_DWIDTH
-
1
:
0
]
}
;
parameter
[
16
*
APB_DWIDTH
-
1
:
0
]
FIXED_PWM_NEGEDGE
=
{
FIXED_PWM_NEGEDGE16
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE15
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE14
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE13
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE12
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE11
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE10
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE9
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE8
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE7
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE6
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE5
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE4
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE3
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE2
[
APB_DWIDTH
-
1
:
0
]
,
FIXED_PWM_NEGEDGE1
[
APB_DWIDTH
-
1
:
0
]
}
;
generate
if
(
CONFIG_MODE
>
0
)
begin
:
CPWMI0
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMII
<=
0
;
end
else
begin
if
(
(
PSEL
==
1
'b
1
)
&&
(
PWRITE
==
1
'b
1
)
&&
(
PENABLE
==
1
'b
1
)
)
begin
case
(
PADDR
[
7
:
2
]
)
37
:
CPWMII
<=
PWDATA
[
3
:
0
]
;
endcase
end
end
end
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMlI
<=
0
;
PWM_STRETCH
<=
0
;
TACHMODE
<=
0
;
end
else
begin
if
(
(
PSEL
==
1
'b
1
)
&&
(
PWRITE
==
1
'b
1
)
&&
(
PENABLE
==
1
'b
1
)
)
begin
case
(
PADDR
[
7
:
2
]
)
36
:
PWM_STRETCH
<=
PWDATA
[
PWM_NUM
-
1
:
0
]
;
39
:
CPWMlI
<=
PWDATA
[
TACH_NUM
-
1
:
0
]
;
40
:
TACHMODE
<=
PWDATA
[
TACH_NUM
-
1
:
0
]
;
endcase
end
end
end
always
@(*)
begin
case
(
CPWMII
)
4
'b
0000
:
CPWMll
=
0
;
4
'b
0001
:
CPWMll
=
1
;
4
'b
0010
:
CPWMll
=
3
;
4
'b
0011
:
CPWMll
=
7
;
4
'b
0100
:
CPWMll
=
15
;
4
'b
0101
:
CPWMll
=
31
;
4
'b
0110
:
CPWMll
=
63
;
4
'b
0111
:
CPWMll
=
127
;
4
'b
1000
:
CPWMll
=
255
;
4
'b
1001
:
CPWMll
=
511
;
4
'b
1010
:
CPWMll
=
1023
;
4
'b
1011
:
CPWMll
=
2047
;
default
:
CPWMll
=
2047
;
endcase
end
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
CPWMOl
<=
0
;
CPWMIl
<=
0
;
tach_cnt_clk
<=
0
;
end
else
begin
if
(
CPWMOl
>=
CPWMIl
)
begin
CPWMOl
<=
0
;
CPWMIl
<=
CPWMll
;
tach_cnt_clk
<=
1
;
end
else
begin
CPWMOl
<=
CPWMOl
+
1
;
tach_cnt_clk
<=
0
;
end
end
end
end
endgenerate
genvar
CPWMl0
;
generate
for
(
CPWMl0
=
0
;
CPWMl0
<=
(
TACH_NUM
-
1
)
;
CPWMl0
=
CPWMl0
+
1
)
begin
:
CPWMO1
always
@
(
negedge
PRESETN
or
posedge
PCLK
)
begin
if
(
!
PRESETN
)
begin
TACHSTATUS
[
CPWMl0
]
<=
0
;
status_clear
[
CPWMl0
]
<=
1
'b
1
;
end
else
begin
if
(
(
PSEL
==
1
'b
1
)
&&
(
PWRITE
==
1
'b
1
)
&&
(
PENABLE
==
1
'b
1
)
&&
(
PADDR
[
7
:
2
]
==
6
'h
26
)
)
begin
if
(
PWDATA
[
CPWMl0
]
==
1
'b
1
)
begin
TACHSTATUS
[
CPWMl0
]
<=
1
'b
0
;
status_clear
[
CPWMl0
]
<=
1
'b
1
;
end
end
else
begin
if
(
update_status
[
CPWMl0
]
==
1
'b
1
)
begin
TACHSTATUS
[
CPWMl0
]
<=
1
'b
1
;
status_clear
[
CPWMl0
]
<=
1
'b
0
;
end
end
end
end
end
endgenerate
generate
if
(
CONFIG_MODE
>
0
)
begin
:
CPWMI1
assign
TACHINT
=
TACHINT_ACT_LEVEL
?
(
CPWMOI
)
:
!
(
CPWMOI
)
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
0
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl1
assign
CPWMl
[
0
]
=
PWM_STRETCH_VALUE1
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
1
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOOI
assign
CPWMl
[
1
]
=
PWM_STRETCH_VALUE2
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
2
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIOI
assign
CPWMl
[
2
]
=
PWM_STRETCH_VALUE3
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
3
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlOI
assign
CPWMl
[
3
]
=
PWM_STRETCH_VALUE4
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
4
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOII
assign
CPWMl
[
4
]
=
PWM_STRETCH_VALUE5
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
5
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIII
assign
CPWMl
[
5
]
=
PWM_STRETCH_VALUE6
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
6
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlII
assign
CPWMl
[
6
]
=
PWM_STRETCH_VALUE7
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
7
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOlI
assign
CPWMl
[
7
]
=
PWM_STRETCH_VALUE8
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
8
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIlI
assign
CPWMl
[
8
]
=
PWM_STRETCH_VALUE9
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
9
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMllI
assign
CPWMl
[
9
]
=
PWM_STRETCH_VALUE10
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
10
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMO0I
assign
CPWMl
[
10
]
=
PWM_STRETCH_VALUE11
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
11
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMI0I
assign
CPWMl
[
11
]
=
PWM_STRETCH_VALUE12
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
12
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl0I
assign
CPWMl
[
12
]
=
PWM_STRETCH_VALUE13
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
13
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMO1I
assign
CPWMl
[
13
]
=
PWM_STRETCH_VALUE14
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
14
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMI1I
assign
CPWMl
[
14
]
=
PWM_STRETCH_VALUE15
;
end
endgenerate
generate
if
(
(
PWM_NUM
>
15
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl1I
assign
CPWMl
[
15
]
=
PWM_STRETCH_VALUE16
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
1
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOOl
assign
TACH_EDGE
=
{
TACH_EDGE1
}
;
assign
CPWMOI
=
(
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
2
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIOl
assign
TACH_EDGE
=
{
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
3
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlOl
assign
TACH_EDGE
=
{
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
4
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOIl
assign
TACH_EDGE
=
{
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
5
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIIl
assign
TACH_EDGE
=
{
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
6
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlIl
assign
TACH_EDGE
=
{
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
7
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOll
assign
TACH_EDGE
=
{
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
8
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIll
assign
TACH_EDGE
=
{
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
9
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlll
assign
TACH_EDGE
=
{
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
10
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMO0l
assign
TACH_EDGE
=
{
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
11
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMI0l
assign
TACH_EDGE
=
{
TACH_EDGE11
,
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
10
]
&
CPWMlI
[
10
]
)
|
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
12
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl0l
assign
TACH_EDGE
=
{
TACH_EDGE12
,
TACH_EDGE11
,
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
11
]
&
CPWMlI
[
11
]
)
|
(
TACHSTATUS
[
10
]
&
CPWMlI
[
10
]
)
|
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
13
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMO1l
assign
TACH_EDGE
=
{
TACH_EDGE13
,
TACH_EDGE12
,
TACH_EDGE11
,
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
12
]
&
CPWMlI
[
12
]
)
|
(
TACHSTATUS
[
11
]
&
CPWMlI
[
11
]
)
|
(
TACHSTATUS
[
10
]
&
CPWMlI
[
10
]
)
|
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
14
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMI1l
assign
TACH_EDGE
=
{
TACH_EDGE14
,
TACH_EDGE13
,
TACH_EDGE12
,
TACH_EDGE11
,
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
13
]
&
CPWMlI
[
13
]
)
|
(
TACHSTATUS
[
12
]
&
CPWMlI
[
12
]
)
|
(
TACHSTATUS
[
11
]
&
CPWMlI
[
11
]
)
|
(
TACHSTATUS
[
10
]
&
CPWMlI
[
10
]
)
|
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
15
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl1l
assign
TACH_EDGE
=
{
TACH_EDGE15
,
TACH_EDGE14
,
TACH_EDGE13
,
TACH_EDGE12
,
TACH_EDGE11
,
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
14
]
&
CPWMlI
[
14
]
)
|
(
TACHSTATUS
[
13
]
&
CPWMlI
[
13
]
)
|
(
TACHSTATUS
[
12
]
&
CPWMlI
[
12
]
)
|
(
TACHSTATUS
[
11
]
&
CPWMlI
[
11
]
)
|
(
TACHSTATUS
[
10
]
&
CPWMlI
[
10
]
)
|
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
16
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOO0
assign
TACH_EDGE
=
{
TACH_EDGE16
,
TACH_EDGE15
,
TACH_EDGE14
,
TACH_EDGE13
,
TACH_EDGE12
,
TACH_EDGE11
,
TACH_EDGE10
,
TACH_EDGE9
,
TACH_EDGE8
,
TACH_EDGE7
,
TACH_EDGE6
,
TACH_EDGE5
,
TACH_EDGE4
,
TACH_EDGE3
,
TACH_EDGE2
,
TACH_EDGE1
}
;
assign
CPWMOI
=
(
(
TACHSTATUS
[
15
]
&
CPWMlI
[
15
]
)
|
(
TACHSTATUS
[
14
]
&
CPWMlI
[
14
]
)
|
(
TACHSTATUS
[
13
]
&
CPWMlI
[
13
]
)
|
(
TACHSTATUS
[
12
]
&
CPWMlI
[
12
]
)
|
(
TACHSTATUS
[
11
]
&
CPWMlI
[
11
]
)
|
(
TACHSTATUS
[
10
]
&
CPWMlI
[
10
]
)
|
(
TACHSTATUS
[
9
]
&
CPWMlI
[
9
]
)
|
(
TACHSTATUS
[
8
]
&
CPWMlI
[
8
]
)
|
(
TACHSTATUS
[
7
]
&
CPWMlI
[
7
]
)
|
(
TACHSTATUS
[
6
]
&
CPWMlI
[
6
]
)
|
(
TACHSTATUS
[
5
]
&
CPWMlI
[
5
]
)
|
(
TACHSTATUS
[
4
]
&
CPWMlI
[
4
]
)
|
(
TACHSTATUS
[
3
]
&
CPWMlI
[
3
]
)
|
(
TACHSTATUS
[
2
]
&
CPWMlI
[
2
]
)
|
(
TACHSTATUS
[
1
]
&
CPWMlI
[
1
]
|
TACHSTATUS
[
0
]
&
CPWMlI
[
0
]
)
)
;
end
endgenerate
generate
if
(
(
TACH_NUM
==
1
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIO0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
2
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlO0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
3
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOI0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
4
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMII0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
5
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMlI0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
6
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOl0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
7
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIl0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
8
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMll0
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
9
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMO00
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
10
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMI00
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
11
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl00
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
6
'h
33
:
CPWMI
=
TACHPULSEDUR
[
10
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
12
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMO10
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
6
'h
33
:
CPWMI
=
TACHPULSEDUR
[
10
]
;
6
'h
34
:
CPWMI
=
TACHPULSEDUR
[
11
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
13
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMI10
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
6
'h
33
:
CPWMI
=
TACHPULSEDUR
[
10
]
;
6
'h
34
:
CPWMI
=
TACHPULSEDUR
[
11
]
;
6
'h
35
:
CPWMI
=
TACHPULSEDUR
[
12
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
14
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMl10
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
6
'h
33
:
CPWMI
=
TACHPULSEDUR
[
10
]
;
6
'h
34
:
CPWMI
=
TACHPULSEDUR
[
11
]
;
6
'h
35
:
CPWMI
=
TACHPULSEDUR
[
12
]
;
6
'h
36
:
CPWMI
=
TACHPULSEDUR
[
13
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
15
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMOO1
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
6
'h
33
:
CPWMI
=
TACHPULSEDUR
[
10
]
;
6
'h
34
:
CPWMI
=
TACHPULSEDUR
[
11
]
;
6
'h
35
:
CPWMI
=
TACHPULSEDUR
[
12
]
;
6
'h
36
:
CPWMI
=
TACHPULSEDUR
[
13
]
;
6
'h
37
:
CPWMI
=
TACHPULSEDUR
[
14
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
(
TACH_NUM
==
16
)
&&
(
CONFIG_MODE
>
0
)
)
begin
:
CPWMIO1
always
@*
begin
case
(
PADDR
[
7
:
2
]
)
6
'h
25
:
CPWMI
=
CPWMII
[
3
:
0
]
;
6
'h
26
:
CPWMI
=
TACHSTATUS
[
TACH_NUM
-
1
:
0
]
;
6
'h
27
:
CPWMI
=
CPWMlI
[
TACH_NUM
-
1
:
0
]
;
6
'h
28
:
CPWMI
=
TACHMODE
[
TACH_NUM
-
1
:
0
]
;
6
'h
29
:
CPWMI
=
TACHPULSEDUR
[
0
]
;
6
'h
2a
:
CPWMI
=
TACHPULSEDUR
[
1
]
;
6
'h
2b
:
CPWMI
=
TACHPULSEDUR
[
2
]
;
6
'h
2c
:
CPWMI
=
TACHPULSEDUR
[
3
]
;
6
'h
2d
:
CPWMI
=
TACHPULSEDUR
[
4
]
;
6
'h
2e
:
CPWMI
=
TACHPULSEDUR
[
5
]
;
6
'h
2f
:
CPWMI
=
TACHPULSEDUR
[
6
]
;
6
'h
30
:
CPWMI
=
TACHPULSEDUR
[
7
]
;
6
'h
31
:
CPWMI
=
TACHPULSEDUR
[
8
]
;
6
'h
32
:
CPWMI
=
TACHPULSEDUR
[
9
]
;
6
'h
33
:
CPWMI
=
TACHPULSEDUR
[
10
]
;
6
'h
34
:
CPWMI
=
TACHPULSEDUR
[
11
]
;
6
'h
35
:
CPWMI
=
TACHPULSEDUR
[
12
]
;
6
'h
36
:
CPWMI
=
TACHPULSEDUR
[
13
]
;
6
'h
37
:
CPWMI
=
TACHPULSEDUR
[
14
]
;
6
'h
38
:
CPWMI
=
TACHPULSEDUR
[
15
]
;
default
:
CPWMI
=
0
;
endcase
end
end
endgenerate
generate
if
(
APB_DWIDTH
==
32
)
begin
assign
PRDATA
=
(
(
PADDR
[
7
:
2
]
<=
6
'h
24
)
||
(
PADDR
[
7
:
2
]
==
6
'h
39
)
)
?
CPWMO0
:
{
16
'b
0
,
CPWMI
[
15
:
0
]
}
;
end
else
if
(
APB_DWIDTH
==
16
)
begin
assign
PRDATA
=
(
(
PADDR
[
7
:
2
]
<=
6
'h
24
)
||
(
PADDR
[
7
:
2
]
==
6
'h
39
)
)
?
CPWMO0
:
CPWMI
[
15
:
0
]
;
end
else
begin
assign
PRDATA
=
CPWMO0
;
end
endgenerate
genvar
CPWMlO1
;
generate
for
(
CPWMlO1
=
1
;
CPWMlO1
<=
(
PWM_NUM
)
;
CPWMlO1
=
CPWMlO1
+
1
)
begin
:
CPWMOI1
if
(
CONFIG_MODE
==
0
)
begin
assign
PWM
[
CPWMlO1
]
=
CPWMO
[
CPWMlO1
]
;
end
else
if
(
CONFIG_MODE
==
1
)
begin
assign
PWM
[
CPWMlO1
]
=
PWM_STRETCH
[
CPWMlO1
-
1
]
?
CPWMl
[
CPWMlO1
-
1
]
:
CPWMO
[
CPWMlO1
]
;
end
end
endgenerate
generate
if
(
CONFIG_MODE
<
2
)
begin
reg_if
#
(
PWM_NUM
,
APB_DWIDTH
,
FIXED_PRESCALE_EN
,
FIXED_PRESCALE
,
FIXED_PERIOD_EN
,
FIXED_PERIOD
,
DAC_MODE
,
SHADOW_REG_EN
,
FIXED_PWM_POS_EN
,
FIXED_PWM_POSEDGE
,
FIXED_PWM_NEG_EN
,
FIXED_PWM_NEGEDGE
)
reg_if
(
.PCLK
(
PCLK
)
,
.PRESETN
(
PRESETN
)
,
.PSEL
(
PSEL
)
,
.PENABLE
(
PENABLE
)
,
.PWRITE
(
PWRITE
)
,
.PADDR
(
PADDR
[
7
:
2
]
)
,
.PWDATA
(
PWDATA
)
,
.PWM_STRETCH
(
PWM_STRETCH
)
,
.CPWMO0
(
CPWMO0
)
,
.pwm_posedge_out_wire
(
pwm_posedge_reg
)
,
.pwm_negedge_out_wire
(
pwm_negedge_reg
)
,
.prescale_out_wire
(
prescale_reg
)
,
.period_out_wire
(
period_reg
)
,
.period_cnt
(
period_cnt
)
,
.pwm_enable_out_wire
(
pwm_enable_reg
)
,
.sync_pulse
(
sync_pulse
)
)
;
end
endgenerate
genvar
CPWMII1
;
generate
if
(
(
CONFIG_MODE
>
0
)
&&
(
APB_DWIDTH
>
15
)
)
for
(
CPWMII1
=
0
;
CPWMII1
<=
(
TACH_NUM
-
1
)
;
CPWMII1
=
CPWMII1
+
1
)
begin
:
CPWMlI1
tach_if
#
(
.TACH_NUM
(
TACH_NUM
)
)
tach_if
(
.PCLK
(
PCLK
)
,
.PRESETN
(
PRESETN
)
,
.TACHSTATUS
(
TACHSTATUS
[
CPWMII1
]
)
,
.TACH_EDGE
(
TACH_EDGE
[
CPWMII1
]
)
,
.TACHIN
(
TACHIN
[
CPWMII1
]
)
,
.TACHMODE
(
TACHMODE
[
CPWMII1
]
)
,
.status_clear
(
status_clear
[
CPWMII1
]
)
,
.tach_cnt_clk
(
tach_cnt_clk
)
,
.TACHPULSEDUR
(
TACHPULSEDUR
[
CPWMII1
]
)
,
.update_status
(
update_status
[
CPWMII1
]
)
)
;
end
endgenerate
assign
PREADY
=
1
'b
1
;
assign
PSLVERR
=
1
'b
0
;
generate
if
(
(
SHADOW_REG_EN
[
PWM_NUM
-
1
:
0
]
==
0
)
&&
(
DAC_MODE
[
PWM_NUM
-
1
:
0
]
==
all_ones
[
PWM_NUM
-
1
:
0
]
)
)
begin
assign
period_cnt
=
0
;
assign
sync_pulse
=
0
;
end
else
begin
if
(
CONFIG_MODE
<
2
)
begin
timebase
#
(
APB_DWIDTH
)
timebase
(
.PCLK
(
PCLK
)
,
.PRESETN
(
PRESETN
)
,
.prescale_reg
(
prescale_reg
)
,
.period_reg
(
period_reg
)
,
.period_cnt
(
period_cnt
)
,
.sync_pulse
(
sync_pulse
)
)
;
end
end
endgenerate
generate
if
(
CONFIG_MODE
<
2
)
begin
pwm_gen
#
(
PWM_NUM
,
APB_DWIDTH
,
DAC_MODE
)
pwm_gen
(
.PCLK
(
PCLK
)
,
.PRESETN
(
PRESETN
)
,
.PWM
(
CPWMO
)
,
.period_cnt
(
period_cnt
)
,
.pwm_enable_reg
(
pwm_enable_reg
)
,
.pwm_posedge_reg
(
pwm_posedge_reg
)
,
.pwm_negedge_reg
(
pwm_negedge_reg
)
,
.sync_pulse
(
sync_pulse
)
)
;
end
endgenerate
endmodule
