`timescale 1 ns/100 ps
// Version: 9.1 SP5 9.1.5.1


module final_top(
       UART_0_TXD,
       UART_0_RXD,
       MSS_RESET_N,
       GPIO_0_BI,
       UART_1_TXD,
       UART_1_RXD,
       RX,
       TX
    );
output UART_0_TXD;
input  UART_0_RXD;
input  MSS_RESET_N;
inout  GPIO_0_BI;
output UART_1_TXD;
input  UART_1_RXD;
input  RX;
output TX;

    wire \CoreAPB3_0_APBmslave0_PADDR_[0] , 
        \CoreAPB3_0_APBmslave0_PADDR_[1] , 
        \CoreAPB3_0_APBmslave0_PADDR_[2] , 
        \CoreAPB3_0_APBmslave0_PADDR_[3] , 
        \CoreAPB3_0_APBmslave0_PADDR_[4] , 
        \CoreAPB3_0_APBmslave0_PADDR_[5] , 
        \CoreAPB3_0_APBmslave0_PADDR_[6] , 
        \CoreAPB3_0_APBmslave0_PADDR_[7] , 
        \CoreAPB3_0_APBmslave0_PADDR_[8] , 
        \CoreAPB3_0_APBmslave0_PADDR_[9] , 
        \CoreAPB3_0_APBmslave0_PADDR_[10] , 
        \CoreAPB3_0_APBmslave0_PADDR_[11] , 
        \CoreAPB3_0_APBmslave0_PADDR_[12] , 
        \CoreAPB3_0_APBmslave0_PADDR_[13] , 
        \CoreAPB3_0_APBmslave0_PADDR_[14] , 
        \CoreAPB3_0_APBmslave0_PADDR_[15] , 
        \CoreAPB3_0_APBmslave0_PADDR_[16] , 
        \CoreAPB3_0_APBmslave0_PADDR_[17] , 
        \CoreAPB3_0_APBmslave0_PADDR_[18] , 
        \CoreAPB3_0_APBmslave0_PADDR_[19] , 
        \CoreAPB3_0_APBmslave0_PADDR_[20] , 
        \CoreAPB3_0_APBmslave0_PADDR_[21] , 
        \CoreAPB3_0_APBmslave0_PADDR_[22] , 
        \CoreAPB3_0_APBmslave0_PADDR_[23] , 
        CoreAPB3_0_APBmslave0_PENABLE, 
        \CoreAPB3_0_APBmslave0_PRDATA_[0] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[7] , 
        CoreAPB3_0_APBmslave0_PREADY, CoreAPB3_0_APBmslave0_PSELx, 
        CoreAPB3_0_APBmslave0_PSLVERR, 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[31] , 
        CoreAPB3_0_APBmslave0_PWRITE, final_mss_0_FAB_CLK_0, 
        final_mss_0_M2F_RESET_N, 
        \final_mss_0_MSS_MASTER_APB_PADDR_[0] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[1] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[2] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[3] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[4] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[5] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[6] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[7] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[8] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[9] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[10] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[11] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[12] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[13] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[14] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[15] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[16] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[17] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[18] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[19] , 
        final_mss_0_MSS_MASTER_APB_PENABLE, 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[0] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[31] , 
        final_mss_0_MSS_MASTER_APB_PREADY, 
        final_mss_0_MSS_MASTER_APB_PSELx, 
        final_mss_0_MSS_MASTER_APB_PSLVERR, 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[0] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[31] , 
        final_mss_0_MSS_MASTER_APB_PWRITE, GND_net, VCC_net;
    
    CoreAPB3 #( .APBSLOT0ENABLE(1), .APBSLOT10ENABLE(0), .APBSLOT11ENABLE(0)
        , .APBSLOT12ENABLE(0), .APBSLOT13ENABLE(0), .APBSLOT14ENABLE(0)
        , .APBSLOT15ENABLE(0), .APBSLOT1ENABLE(0), .APBSLOT2ENABLE(0)
        , .APBSLOT3ENABLE(0), .APBSLOT4ENABLE(0), .APBSLOT5ENABLE(0), .APBSLOT6ENABLE(0)
        , .APBSLOT7ENABLE(0), .APBSLOT8ENABLE(0), .APBSLOT9ENABLE(0), .APB_DWIDTH(32)
        , .IADDR_ENABLE(0), .RANGESIZE(256) )  CoreAPB3_0 (.PRESETN(
        GND_net), .PCLK(GND_net), .PADDR({GND_net, GND_net, GND_net, 
        GND_net, \final_mss_0_MSS_MASTER_APB_PADDR_[19] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[18] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[17] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[16] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[15] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[14] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[13] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[12] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[11] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[10] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[9] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[8] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[7] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[6] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[5] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[4] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[3] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[2] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[1] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[0] }), .PWRITE(
        final_mss_0_MSS_MASTER_APB_PWRITE), .PENABLE(
        final_mss_0_MSS_MASTER_APB_PENABLE), .PWDATA({
        \final_mss_0_MSS_MASTER_APB_PWDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[0] }), .PRDATA({
        \final_mss_0_MSS_MASTER_APB_PRDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[0] }), .PSEL(
        final_mss_0_MSS_MASTER_APB_PSELx), .PREADY(
        final_mss_0_MSS_MASTER_APB_PREADY), .PSLVERR(
        final_mss_0_MSS_MASTER_APB_PSLVERR), .PADDRS({nc0, nc1, nc2, 
        nc3, nc4, nc5, nc6, nc7, nc8, nc9, nc10, nc11, nc12, nc13, 
        nc14, nc15, nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23}), 
        .PADDRS0({\CoreAPB3_0_APBmslave0_PADDR_[23] , 
        \CoreAPB3_0_APBmslave0_PADDR_[22] , 
        \CoreAPB3_0_APBmslave0_PADDR_[21] , 
        \CoreAPB3_0_APBmslave0_PADDR_[20] , 
        \CoreAPB3_0_APBmslave0_PADDR_[19] , 
        \CoreAPB3_0_APBmslave0_PADDR_[18] , 
        \CoreAPB3_0_APBmslave0_PADDR_[17] , 
        \CoreAPB3_0_APBmslave0_PADDR_[16] , 
        \CoreAPB3_0_APBmslave0_PADDR_[15] , 
        \CoreAPB3_0_APBmslave0_PADDR_[14] , 
        \CoreAPB3_0_APBmslave0_PADDR_[13] , 
        \CoreAPB3_0_APBmslave0_PADDR_[12] , 
        \CoreAPB3_0_APBmslave0_PADDR_[11] , 
        \CoreAPB3_0_APBmslave0_PADDR_[10] , 
        \CoreAPB3_0_APBmslave0_PADDR_[9] , 
        \CoreAPB3_0_APBmslave0_PADDR_[8] , 
        \CoreAPB3_0_APBmslave0_PADDR_[7] , 
        \CoreAPB3_0_APBmslave0_PADDR_[6] , 
        \CoreAPB3_0_APBmslave0_PADDR_[5] , 
        \CoreAPB3_0_APBmslave0_PADDR_[4] , 
        \CoreAPB3_0_APBmslave0_PADDR_[3] , 
        \CoreAPB3_0_APBmslave0_PADDR_[2] , 
        \CoreAPB3_0_APBmslave0_PADDR_[1] , 
        \CoreAPB3_0_APBmslave0_PADDR_[0] }), .PWRITES(
        CoreAPB3_0_APBmslave0_PWRITE), .PENABLES(
        CoreAPB3_0_APBmslave0_PENABLE), .PWDATAS({
        \CoreAPB3_0_APBmslave0_PWDATA_[31] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] }), .PSELS0(
        CoreAPB3_0_APBmslave0_PSELx), .PRDATAS0({GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, \CoreAPB3_0_APBmslave0_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[0] }), .PREADYS0(
        CoreAPB3_0_APBmslave0_PREADY), .PSLVERRS0(
        CoreAPB3_0_APBmslave0_PSLVERR), .PSELS1(), .PRDATAS1({GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net}), .PREADYS1(VCC_net), .PSLVERRS1(
        GND_net), .PSELS2(), .PRDATAS2({GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net}), .PREADYS2(VCC_net), .PSLVERRS2(GND_net), .PSELS3(), 
        .PRDATAS3({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS3(VCC_net), .PSLVERRS3(GND_net), .PSELS4(), .PRDATAS4({
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net}), .PREADYS4(VCC_net), 
        .PSLVERRS4(GND_net), .PSELS5(), .PRDATAS5({GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net}), .PREADYS5(VCC_net), .PSLVERRS5(GND_net), 
        .PSELS6(), .PRDATAS6({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net})
        , .PREADYS6(VCC_net), .PSLVERRS6(GND_net), .PSELS7(), 
        .PRDATAS7({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS7(VCC_net), .PSLVERRS7(GND_net), .PSELS8(), .PRDATAS8({
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net}), .PREADYS8(VCC_net), 
        .PSLVERRS8(GND_net), .PSELS9(), .PRDATAS9({GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net}), .PREADYS9(VCC_net), .PSLVERRS9(GND_net), 
        .PSELS10(), .PRDATAS10({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net})
        , .PREADYS10(VCC_net), .PSLVERRS10(GND_net), .PSELS11(), 
        .PRDATAS11({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS11(VCC_net), .PSLVERRS11(GND_net), .PSELS12(), 
        .PRDATAS12({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS12(VCC_net), .PSLVERRS12(GND_net), .PSELS13(), 
        .PRDATAS13({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS13(VCC_net), .PSLVERRS13(GND_net), .PSELS14(), 
        .PRDATAS14({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS14(VCC_net), .PSLVERRS14(GND_net), .PSELS15(), 
        .PRDATAS15({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PREADYS15(VCC_net), .PSLVERRS15(GND_net));
    VCC VCC (.Y(VCC_net));
    GND GND (.Y(GND_net));
    final_mss final_mss_0 (.MSS_RESET_N(MSS_RESET_N), .M2F_RESET_N(
        final_mss_0_M2F_RESET_N), .GPIO_0_BI(GPIO_0_BI), .UART_0_TXD(
        UART_0_TXD), .UART_0_RXD(UART_0_RXD), .UART_1_TXD(UART_1_TXD), 
        .UART_1_RXD(UART_1_RXD), .MSSPSEL(
        final_mss_0_MSS_MASTER_APB_PSELx), .MSSPENABLE(
        final_mss_0_MSS_MASTER_APB_PENABLE), .MSSPWRITE(
        final_mss_0_MSS_MASTER_APB_PWRITE), .MSSPREADY(
        final_mss_0_MSS_MASTER_APB_PREADY), .MSSPSLVERR(
        final_mss_0_MSS_MASTER_APB_PSLVERR), .FAB_CLK(
        final_mss_0_FAB_CLK_0), .MSSPADDR({
        \final_mss_0_MSS_MASTER_APB_PADDR_[19] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[18] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[17] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[16] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[15] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[14] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[13] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[12] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[11] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[10] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[9] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[8] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[7] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[6] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[5] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[4] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[3] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[2] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[1] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[0] }), .MSSPRDATA({
        \final_mss_0_MSS_MASTER_APB_PRDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[0] }), .MSSPWDATA({
        \final_mss_0_MSS_MASTER_APB_PWDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[0] }));
    final_top_CoreUARTapb_0_CoreUARTapb #( .BAUD_VALUE(4800), .BAUD_VAL_FRCTN(0)
        , .BAUD_VAL_FRCTN_EN(0), .FAMILY(18), .FIXEDMODE(1), .PRG_BIT8(1)
        , .PRG_PARITY(0), .RX_FIFO(1), .RX_LEGACY_MODE(0), .TX_FIFO(1)
         )  CoreUARTapb_0 (.PCLK(final_mss_0_FAB_CLK_0), .PRESETN(
        final_mss_0_M2F_RESET_N), .PADDR({
        \CoreAPB3_0_APBmslave0_PADDR_[4] , 
        \CoreAPB3_0_APBmslave0_PADDR_[3] , 
        \CoreAPB3_0_APBmslave0_PADDR_[2] , 
        \CoreAPB3_0_APBmslave0_PADDR_[1] , 
        \CoreAPB3_0_APBmslave0_PADDR_[0] }), .PSEL(
        CoreAPB3_0_APBmslave0_PSELx), .PENABLE(
        CoreAPB3_0_APBmslave0_PENABLE), .PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] }), .PRDATA({
        \CoreAPB3_0_APBmslave0_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[0] }), .TXRDY(), .RXRDY(), 
        .PARITY_ERR(), .OVERFLOW(), .RX(RX), .TX(TX), .PREADY(
        CoreAPB3_0_APBmslave0_PREADY), .PSLVERR(
        CoreAPB3_0_APBmslave0_PSLVERR), .FRAMING_ERR());
    
endmodule
