`timescale 1 ns/100 ps
// Version: 9.1 SP5 9.1.5.1


module final_top(
       MSS_RESET_N,
       UART_0_TXD,
       UART_0_RXD,
       ADCDirectInput_0,
       VAREF1,
       UART_1_TXD,
       UART_1_RXD,
       RX,
       TX,
       PWM,
       TACHIN,
       GPIO_15_OUT,
       PWM_0
    );
input  MSS_RESET_N;
output UART_0_TXD;
input  UART_0_RXD;
input  ADCDirectInput_0;
input  VAREF1;
output UART_1_TXD;
input  UART_1_RXD;
input  RX;
output TX;
output [8:1] PWM;
input  [1:1] TACHIN;
output GPIO_15_OUT;
output [2:1] PWM_0;

    wire \CoreAPB3_0_APBmslave0_PADDR_[0] , 
        \CoreAPB3_0_APBmslave0_PADDR_[1] , 
        \CoreAPB3_0_APBmslave0_PADDR_[2] , 
        \CoreAPB3_0_APBmslave0_PADDR_[3] , 
        \CoreAPB3_0_APBmslave0_PADDR_[4] , 
        \CoreAPB3_0_APBmslave0_PADDR_[5] , 
        \CoreAPB3_0_APBmslave0_PADDR_[6] , 
        \CoreAPB3_0_APBmslave0_PADDR_[7] , 
        \CoreAPB3_0_APBmslave0_PADDR_[8] , 
        \CoreAPB3_0_APBmslave0_PADDR_[9] , 
        \CoreAPB3_0_APBmslave0_PADDR_[10] , 
        \CoreAPB3_0_APBmslave0_PADDR_[11] , 
        \CoreAPB3_0_APBmslave0_PADDR_[12] , 
        \CoreAPB3_0_APBmslave0_PADDR_[13] , 
        \CoreAPB3_0_APBmslave0_PADDR_[14] , 
        \CoreAPB3_0_APBmslave0_PADDR_[15] , 
        \CoreAPB3_0_APBmslave0_PADDR_[16] , 
        \CoreAPB3_0_APBmslave0_PADDR_[17] , 
        \CoreAPB3_0_APBmslave0_PADDR_[18] , 
        \CoreAPB3_0_APBmslave0_PADDR_[19] , 
        \CoreAPB3_0_APBmslave0_PADDR_[20] , 
        \CoreAPB3_0_APBmslave0_PADDR_[21] , 
        \CoreAPB3_0_APBmslave0_PADDR_[22] , 
        \CoreAPB3_0_APBmslave0_PADDR_[23] , 
        CoreAPB3_0_APBmslave0_PENABLE, 
        \CoreAPB3_0_APBmslave0_PRDATA_[0] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[31] , 
        CoreAPB3_0_APBmslave0_PREADY, CoreAPB3_0_APBmslave0_PSELx, 
        CoreAPB3_0_APBmslave0_PSLVERR, 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[31] , 
        CoreAPB3_0_APBmslave0_PWRITE, 
        \CoreAPB3_0_APBmslave1_PADDR_[0] , 
        \CoreAPB3_0_APBmslave1_PADDR_[1] , 
        \CoreAPB3_0_APBmslave1_PADDR_[2] , 
        \CoreAPB3_0_APBmslave1_PADDR_[3] , 
        \CoreAPB3_0_APBmslave1_PADDR_[4] , 
        \CoreAPB3_0_APBmslave1_PADDR_[5] , 
        \CoreAPB3_0_APBmslave1_PADDR_[6] , 
        \CoreAPB3_0_APBmslave1_PADDR_[7] , 
        \CoreAPB3_0_APBmslave1_PADDR_[8] , 
        \CoreAPB3_0_APBmslave1_PADDR_[9] , 
        \CoreAPB3_0_APBmslave1_PADDR_[10] , 
        \CoreAPB3_0_APBmslave1_PADDR_[11] , 
        \CoreAPB3_0_APBmslave1_PADDR_[12] , 
        \CoreAPB3_0_APBmslave1_PADDR_[13] , 
        \CoreAPB3_0_APBmslave1_PADDR_[14] , 
        \CoreAPB3_0_APBmslave1_PADDR_[15] , 
        \CoreAPB3_0_APBmslave1_PADDR_[16] , 
        \CoreAPB3_0_APBmslave1_PADDR_[17] , 
        \CoreAPB3_0_APBmslave1_PADDR_[18] , 
        \CoreAPB3_0_APBmslave1_PADDR_[19] , 
        \CoreAPB3_0_APBmslave1_PADDR_[20] , 
        \CoreAPB3_0_APBmslave1_PADDR_[21] , 
        \CoreAPB3_0_APBmslave1_PADDR_[22] , 
        \CoreAPB3_0_APBmslave1_PADDR_[23] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[0] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[8] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[9] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[10] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[11] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[12] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[13] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[14] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[15] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[16] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[17] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[18] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[19] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[20] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[21] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[22] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[23] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[24] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[25] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[26] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[27] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[28] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[29] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[30] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[31] , 
        CoreAPB3_0_APBmslave1_PREADY, CoreAPB3_0_APBmslave1_PSELx, 
        CoreAPB3_0_APBmslave1_PSLVERR, 
        \CoreAPB3_0_APBmslave2_PRDATA_[0] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[7] , 
        CoreAPB3_0_APBmslave2_PREADY, CoreAPB3_0_APBmslave2_PSELx, 
        CoreAPB3_0_APBmslave2_PSLVERR, final_mss_0_FAB_CLK, 
        final_mss_0_M2F_RESET_N, 
        \final_mss_0_MSS_MASTER_APB_PADDR_[0] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[1] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[2] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[3] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[4] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[5] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[6] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[7] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[8] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[9] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[10] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[11] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[12] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[13] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[14] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[15] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[16] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[17] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[18] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[19] , 
        final_mss_0_MSS_MASTER_APB_PENABLE, 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[0] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[31] , 
        final_mss_0_MSS_MASTER_APB_PREADY, 
        final_mss_0_MSS_MASTER_APB_PSELx, 
        final_mss_0_MSS_MASTER_APB_PSLVERR, 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[0] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[31] , 
        final_mss_0_MSS_MASTER_APB_PWRITE, GND_net, VCC_net;
    
    CoreAPB3 #( .APBSLOT0ENABLE(1), .APBSLOT10ENABLE(0), .APBSLOT11ENABLE(0)
        , .APBSLOT12ENABLE(0), .APBSLOT13ENABLE(0), .APBSLOT14ENABLE(0)
        , .APBSLOT15ENABLE(0), .APBSLOT1ENABLE(1), .APBSLOT2ENABLE(1)
        , .APBSLOT3ENABLE(0), .APBSLOT4ENABLE(0), .APBSLOT5ENABLE(0), .APBSLOT6ENABLE(0)
        , .APBSLOT7ENABLE(0), .APBSLOT8ENABLE(0), .APBSLOT9ENABLE(0), .APB_DWIDTH(32)
        , .IADDR_ENABLE(0), .RANGESIZE(256) )  CoreAPB3_0 (.PRESETN(
        GND_net), .PCLK(GND_net), .PWRITE(
        final_mss_0_MSS_MASTER_APB_PWRITE), .PENABLE(
        final_mss_0_MSS_MASTER_APB_PENABLE), .PSEL(
        final_mss_0_MSS_MASTER_APB_PSELx), .PREADY(
        final_mss_0_MSS_MASTER_APB_PREADY), .PSLVERR(
        final_mss_0_MSS_MASTER_APB_PSLVERR), .PWRITES(
        CoreAPB3_0_APBmslave0_PWRITE), .PENABLES(
        CoreAPB3_0_APBmslave0_PENABLE), .PSELS0(
        CoreAPB3_0_APBmslave0_PSELx), .PREADYS0(
        CoreAPB3_0_APBmslave0_PREADY), .PSLVERRS0(
        CoreAPB3_0_APBmslave0_PSLVERR), .PSELS1(
        CoreAPB3_0_APBmslave1_PSELx), .PREADYS1(
        CoreAPB3_0_APBmslave1_PREADY), .PSLVERRS1(
        CoreAPB3_0_APBmslave1_PSLVERR), .PSELS2(
        CoreAPB3_0_APBmslave2_PSELx), .PREADYS2(
        CoreAPB3_0_APBmslave2_PREADY), .PSLVERRS2(
        CoreAPB3_0_APBmslave2_PSLVERR), .PSELS3(), .PREADYS3(VCC_net), 
        .PSLVERRS3(GND_net), .PSELS4(), .PREADYS4(VCC_net), .PSLVERRS4(
        GND_net), .PSELS5(), .PREADYS5(VCC_net), .PSLVERRS5(GND_net), 
        .PSELS6(), .PREADYS6(VCC_net), .PSLVERRS6(GND_net), .PSELS7(), 
        .PREADYS7(VCC_net), .PSLVERRS7(GND_net), .PSELS8(), .PREADYS8(
        VCC_net), .PSLVERRS8(GND_net), .PSELS9(), .PREADYS9(VCC_net), 
        .PSLVERRS9(GND_net), .PSELS10(), .PREADYS10(VCC_net), 
        .PSLVERRS10(GND_net), .PSELS11(), .PREADYS11(VCC_net), 
        .PSLVERRS11(GND_net), .PSELS12(), .PREADYS12(VCC_net), 
        .PSLVERRS12(GND_net), .PSELS13(), .PREADYS13(VCC_net), 
        .PSLVERRS13(GND_net), .PSELS14(), .PREADYS14(VCC_net), 
        .PSLVERRS14(GND_net), .PSELS15(), .PREADYS15(VCC_net), 
        .PSLVERRS15(GND_net), .PADDR({GND_net, GND_net, GND_net, 
        GND_net, \final_mss_0_MSS_MASTER_APB_PADDR_[19] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[18] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[17] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[16] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[15] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[14] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[13] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[12] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[11] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[10] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[9] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[8] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[7] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[6] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[5] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[4] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[3] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[2] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[1] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[0] }), .PWDATA({
        \final_mss_0_MSS_MASTER_APB_PWDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[0] }), .PRDATA({
        \final_mss_0_MSS_MASTER_APB_PRDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[0] }), .PADDRS({
        \CoreAPB3_0_APBmslave1_PADDR_[23] , 
        \CoreAPB3_0_APBmslave1_PADDR_[22] , 
        \CoreAPB3_0_APBmslave1_PADDR_[21] , 
        \CoreAPB3_0_APBmslave1_PADDR_[20] , 
        \CoreAPB3_0_APBmslave1_PADDR_[19] , 
        \CoreAPB3_0_APBmslave1_PADDR_[18] , 
        \CoreAPB3_0_APBmslave1_PADDR_[17] , 
        \CoreAPB3_0_APBmslave1_PADDR_[16] , 
        \CoreAPB3_0_APBmslave1_PADDR_[15] , 
        \CoreAPB3_0_APBmslave1_PADDR_[14] , 
        \CoreAPB3_0_APBmslave1_PADDR_[13] , 
        \CoreAPB3_0_APBmslave1_PADDR_[12] , 
        \CoreAPB3_0_APBmslave1_PADDR_[11] , 
        \CoreAPB3_0_APBmslave1_PADDR_[10] , 
        \CoreAPB3_0_APBmslave1_PADDR_[9] , 
        \CoreAPB3_0_APBmslave1_PADDR_[8] , 
        \CoreAPB3_0_APBmslave1_PADDR_[7] , 
        \CoreAPB3_0_APBmslave1_PADDR_[6] , 
        \CoreAPB3_0_APBmslave1_PADDR_[5] , 
        \CoreAPB3_0_APBmslave1_PADDR_[4] , 
        \CoreAPB3_0_APBmslave1_PADDR_[3] , 
        \CoreAPB3_0_APBmslave1_PADDR_[2] , 
        \CoreAPB3_0_APBmslave1_PADDR_[1] , 
        \CoreAPB3_0_APBmslave1_PADDR_[0] }), .PADDRS0({
        \CoreAPB3_0_APBmslave0_PADDR_[23] , 
        \CoreAPB3_0_APBmslave0_PADDR_[22] , 
        \CoreAPB3_0_APBmslave0_PADDR_[21] , 
        \CoreAPB3_0_APBmslave0_PADDR_[20] , 
        \CoreAPB3_0_APBmslave0_PADDR_[19] , 
        \CoreAPB3_0_APBmslave0_PADDR_[18] , 
        \CoreAPB3_0_APBmslave0_PADDR_[17] , 
        \CoreAPB3_0_APBmslave0_PADDR_[16] , 
        \CoreAPB3_0_APBmslave0_PADDR_[15] , 
        \CoreAPB3_0_APBmslave0_PADDR_[14] , 
        \CoreAPB3_0_APBmslave0_PADDR_[13] , 
        \CoreAPB3_0_APBmslave0_PADDR_[12] , 
        \CoreAPB3_0_APBmslave0_PADDR_[11] , 
        \CoreAPB3_0_APBmslave0_PADDR_[10] , 
        \CoreAPB3_0_APBmslave0_PADDR_[9] , 
        \CoreAPB3_0_APBmslave0_PADDR_[8] , 
        \CoreAPB3_0_APBmslave0_PADDR_[7] , 
        \CoreAPB3_0_APBmslave0_PADDR_[6] , 
        \CoreAPB3_0_APBmslave0_PADDR_[5] , 
        \CoreAPB3_0_APBmslave0_PADDR_[4] , 
        \CoreAPB3_0_APBmslave0_PADDR_[3] , 
        \CoreAPB3_0_APBmslave0_PADDR_[2] , 
        \CoreAPB3_0_APBmslave0_PADDR_[1] , 
        \CoreAPB3_0_APBmslave0_PADDR_[0] }), .PWDATAS({
        \CoreAPB3_0_APBmslave0_PWDATA_[31] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] }), .PRDATAS0({
        \CoreAPB3_0_APBmslave0_PRDATA_[31] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[0] }), .PRDATAS1({
        \CoreAPB3_0_APBmslave1_PRDATA_[31] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[30] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[29] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[28] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[27] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[26] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[25] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[24] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[23] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[22] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[21] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[20] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[19] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[18] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[17] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[16] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[15] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[14] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[13] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[12] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[11] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[10] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[9] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[8] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[0] }), .PRDATAS2({GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, \CoreAPB3_0_APBmslave2_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[0] }), .PRDATAS3({GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net}), .PRDATAS4({GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net}), .PRDATAS5({GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net}), .PRDATAS6({GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net})
        , .PRDATAS7({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS8({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS9({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS10({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS11({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS12({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS13({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS14({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}), 
        .PRDATAS15({GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, GND_net, 
        GND_net, GND_net, GND_net, GND_net, GND_net, GND_net}));
    VCC VCC (.Y(VCC_net));
    corepwm #( .APB_DWIDTH(32), .CONFIG_MODE(0), .DAC_MODE1(0), .DAC_MODE10(0)
        , .DAC_MODE11(0), .DAC_MODE12(0), .DAC_MODE13(0), .DAC_MODE14(0)
        , .DAC_MODE15(0), .DAC_MODE16(0), .DAC_MODE2(0), .DAC_MODE3(0)
        , .DAC_MODE4(0), .DAC_MODE5(0), .DAC_MODE6(0), .DAC_MODE7(0), .DAC_MODE8(0)
        , .DAC_MODE9(0), .FAMILY(15), .FIXED_PERIOD(1), .FIXED_PERIOD_EN(0)
        , .FIXED_PRESCALE(0), .FIXED_PRESCALE_EN(0), .FIXED_PWM_NEGEDGE1(0)
        , .FIXED_PWM_NEGEDGE10(0), .FIXED_PWM_NEGEDGE11(0), .FIXED_PWM_NEGEDGE12(0)
        , .FIXED_PWM_NEGEDGE13(0), .FIXED_PWM_NEGEDGE14(0), .FIXED_PWM_NEGEDGE15(0)
        , .FIXED_PWM_NEGEDGE16(0), .FIXED_PWM_NEGEDGE2(0), .FIXED_PWM_NEGEDGE3(0)
        , .FIXED_PWM_NEGEDGE4(0), .FIXED_PWM_NEGEDGE5(0), .FIXED_PWM_NEGEDGE6(0)
        , .FIXED_PWM_NEGEDGE7(0), .FIXED_PWM_NEGEDGE8(0), .FIXED_PWM_NEGEDGE9(0)
        , .FIXED_PWM_NEG_EN1(0), .FIXED_PWM_NEG_EN10(0), .FIXED_PWM_NEG_EN11(0)
        , .FIXED_PWM_NEG_EN12(0), .FIXED_PWM_NEG_EN13(0), .FIXED_PWM_NEG_EN14(0)
        , .FIXED_PWM_NEG_EN15(0), .FIXED_PWM_NEG_EN16(0), .FIXED_PWM_NEG_EN2(0)
        , .FIXED_PWM_NEG_EN3(0), .FIXED_PWM_NEG_EN4(0), .FIXED_PWM_NEG_EN5(0)
        , .FIXED_PWM_NEG_EN6(0), .FIXED_PWM_NEG_EN7(0), .FIXED_PWM_NEG_EN8(0)
        , .FIXED_PWM_NEG_EN9(0), .FIXED_PWM_POSEDGE1(0), .FIXED_PWM_POSEDGE10(0)
        , .FIXED_PWM_POSEDGE11(0), .FIXED_PWM_POSEDGE12(0), .FIXED_PWM_POSEDGE13(0)
        , .FIXED_PWM_POSEDGE14(0), .FIXED_PWM_POSEDGE15(0), .FIXED_PWM_POSEDGE16(0)
        , .FIXED_PWM_POSEDGE2(0), .FIXED_PWM_POSEDGE3(0), .FIXED_PWM_POSEDGE4(0)
        , .FIXED_PWM_POSEDGE5(0), .FIXED_PWM_POSEDGE6(0), .FIXED_PWM_POSEDGE7(0)
        , .FIXED_PWM_POSEDGE8(0), .FIXED_PWM_POSEDGE9(0), .FIXED_PWM_POS_EN1(1)
        , .FIXED_PWM_POS_EN10(1), .FIXED_PWM_POS_EN11(1), .FIXED_PWM_POS_EN12(1)
        , .FIXED_PWM_POS_EN13(1), .FIXED_PWM_POS_EN14(1), .FIXED_PWM_POS_EN15(1)
        , .FIXED_PWM_POS_EN16(1), .FIXED_PWM_POS_EN2(1), .FIXED_PWM_POS_EN3(1)
        , .FIXED_PWM_POS_EN4(1), .FIXED_PWM_POS_EN5(1), .FIXED_PWM_POS_EN6(1)
        , .FIXED_PWM_POS_EN7(1), .FIXED_PWM_POS_EN8(1), .FIXED_PWM_POS_EN9(1)
        , .PWM_NUM(2), .PWM_STRETCH_VALUE1(0), .PWM_STRETCH_VALUE10(0)
        , .PWM_STRETCH_VALUE11(0), .PWM_STRETCH_VALUE12(0), .PWM_STRETCH_VALUE13(0)
        , .PWM_STRETCH_VALUE14(0), .PWM_STRETCH_VALUE15(0), .PWM_STRETCH_VALUE16(0)
        , .PWM_STRETCH_VALUE2(0), .PWM_STRETCH_VALUE3(0), .PWM_STRETCH_VALUE4(0)
        , .PWM_STRETCH_VALUE5(0), .PWM_STRETCH_VALUE6(0), .PWM_STRETCH_VALUE7(0)
        , .PWM_STRETCH_VALUE8(0), .PWM_STRETCH_VALUE9(0), .SHADOW_REG_EN1(0)
        , .SHADOW_REG_EN10(0), .SHADOW_REG_EN11(0), .SHADOW_REG_EN12(0)
        , .SHADOW_REG_EN13(0), .SHADOW_REG_EN14(0), .SHADOW_REG_EN15(0)
        , .SHADOW_REG_EN16(0), .SHADOW_REG_EN2(0), .SHADOW_REG_EN3(0)
        , .SHADOW_REG_EN4(0), .SHADOW_REG_EN5(0), .SHADOW_REG_EN6(0), .SHADOW_REG_EN7(0)
        , .SHADOW_REG_EN8(0), .SHADOW_REG_EN9(0), .TACHINT_ACT_LEVEL(0)
        , .TACH_EDGE1(0), .TACH_EDGE10(0), .TACH_EDGE11(0), .TACH_EDGE12(0)
        , .TACH_EDGE13(0), .TACH_EDGE14(0), .TACH_EDGE15(0), .TACH_EDGE16(0)
        , .TACH_EDGE2(0), .TACH_EDGE3(0), .TACH_EDGE4(0), .TACH_EDGE5(0)
        , .TACH_EDGE6(0), .TACH_EDGE7(0), .TACH_EDGE8(0), .TACH_EDGE9(0)
        , .TACH_NUM(1) )  corepwm_1 (.PADDR({
        \CoreAPB3_0_APBmslave1_PADDR_[7] , 
        \CoreAPB3_0_APBmslave1_PADDR_[6] , 
        \CoreAPB3_0_APBmslave1_PADDR_[5] , 
        \CoreAPB3_0_APBmslave1_PADDR_[4] , 
        \CoreAPB3_0_APBmslave1_PADDR_[3] , 
        \CoreAPB3_0_APBmslave1_PADDR_[2] , 
        \CoreAPB3_0_APBmslave1_PADDR_[1] , 
        \CoreAPB3_0_APBmslave1_PADDR_[0] }), .PCLK(final_mss_0_FAB_CLK)
        , .PENABLE(CoreAPB3_0_APBmslave0_PENABLE), .PRDATA({
        \CoreAPB3_0_APBmslave1_PRDATA_[31] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[30] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[29] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[28] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[27] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[26] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[25] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[24] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[23] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[22] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[21] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[20] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[19] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[18] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[17] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[16] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[15] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[14] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[13] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[12] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[11] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[10] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[9] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[8] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave1_PRDATA_[0] }), .PRESETN(
        final_mss_0_M2F_RESET_N), .PSEL(CoreAPB3_0_APBmslave1_PSELx), 
        .PWDATA({\CoreAPB3_0_APBmslave0_PWDATA_[31] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] }), .PREADY(
        CoreAPB3_0_APBmslave1_PREADY), .PSLVERR(
        CoreAPB3_0_APBmslave1_PSLVERR), .TACHINT(), .TACHIN({TACHIN[1]})
        , .PWM({PWM_0[2], PWM_0[1]}), .PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE));
    corepwm #( .APB_DWIDTH(32), .CONFIG_MODE(0), .DAC_MODE1(0), .DAC_MODE10(0)
        , .DAC_MODE11(0), .DAC_MODE12(0), .DAC_MODE13(0), .DAC_MODE14(0)
        , .DAC_MODE15(0), .DAC_MODE16(0), .DAC_MODE2(0), .DAC_MODE3(0)
        , .DAC_MODE4(0), .DAC_MODE5(0), .DAC_MODE6(0), .DAC_MODE7(0), .DAC_MODE8(0)
        , .DAC_MODE9(0), .FAMILY(15), .FIXED_PERIOD(1), .FIXED_PERIOD_EN(0)
        , .FIXED_PRESCALE(0), .FIXED_PRESCALE_EN(1), .FIXED_PWM_NEGEDGE1(0)
        , .FIXED_PWM_NEGEDGE10(0), .FIXED_PWM_NEGEDGE11(0), .FIXED_PWM_NEGEDGE12(0)
        , .FIXED_PWM_NEGEDGE13(0), .FIXED_PWM_NEGEDGE14(0), .FIXED_PWM_NEGEDGE15(0)
        , .FIXED_PWM_NEGEDGE16(0), .FIXED_PWM_NEGEDGE2(0), .FIXED_PWM_NEGEDGE3(0)
        , .FIXED_PWM_NEGEDGE4(0), .FIXED_PWM_NEGEDGE5(0), .FIXED_PWM_NEGEDGE6(0)
        , .FIXED_PWM_NEGEDGE7(0), .FIXED_PWM_NEGEDGE8(0), .FIXED_PWM_NEGEDGE9(0)
        , .FIXED_PWM_NEG_EN1(0), .FIXED_PWM_NEG_EN10(0), .FIXED_PWM_NEG_EN11(0)
        , .FIXED_PWM_NEG_EN12(0), .FIXED_PWM_NEG_EN13(0), .FIXED_PWM_NEG_EN14(0)
        , .FIXED_PWM_NEG_EN15(0), .FIXED_PWM_NEG_EN16(0), .FIXED_PWM_NEG_EN2(0)
        , .FIXED_PWM_NEG_EN3(0), .FIXED_PWM_NEG_EN4(0), .FIXED_PWM_NEG_EN5(0)
        , .FIXED_PWM_NEG_EN6(0), .FIXED_PWM_NEG_EN7(0), .FIXED_PWM_NEG_EN8(0)
        , .FIXED_PWM_NEG_EN9(0), .FIXED_PWM_POSEDGE1(0), .FIXED_PWM_POSEDGE10(0)
        , .FIXED_PWM_POSEDGE11(0), .FIXED_PWM_POSEDGE12(0), .FIXED_PWM_POSEDGE13(0)
        , .FIXED_PWM_POSEDGE14(0), .FIXED_PWM_POSEDGE15(0), .FIXED_PWM_POSEDGE16(0)
        , .FIXED_PWM_POSEDGE2(0), .FIXED_PWM_POSEDGE3(0), .FIXED_PWM_POSEDGE4(0)
        , .FIXED_PWM_POSEDGE5(0), .FIXED_PWM_POSEDGE6(0), .FIXED_PWM_POSEDGE7(0)
        , .FIXED_PWM_POSEDGE8(0), .FIXED_PWM_POSEDGE9(0), .FIXED_PWM_POS_EN1(1)
        , .FIXED_PWM_POS_EN10(1), .FIXED_PWM_POS_EN11(1), .FIXED_PWM_POS_EN12(1)
        , .FIXED_PWM_POS_EN13(1), .FIXED_PWM_POS_EN14(1), .FIXED_PWM_POS_EN15(1)
        , .FIXED_PWM_POS_EN16(1), .FIXED_PWM_POS_EN2(1), .FIXED_PWM_POS_EN3(1)
        , .FIXED_PWM_POS_EN4(1), .FIXED_PWM_POS_EN5(1), .FIXED_PWM_POS_EN6(1)
        , .FIXED_PWM_POS_EN7(1), .FIXED_PWM_POS_EN8(1), .FIXED_PWM_POS_EN9(1)
        , .PWM_NUM(8), .PWM_STRETCH_VALUE1(0), .PWM_STRETCH_VALUE10(0)
        , .PWM_STRETCH_VALUE11(0), .PWM_STRETCH_VALUE12(0), .PWM_STRETCH_VALUE13(0)
        , .PWM_STRETCH_VALUE14(0), .PWM_STRETCH_VALUE15(0), .PWM_STRETCH_VALUE16(0)
        , .PWM_STRETCH_VALUE2(0), .PWM_STRETCH_VALUE3(0), .PWM_STRETCH_VALUE4(0)
        , .PWM_STRETCH_VALUE5(0), .PWM_STRETCH_VALUE6(0), .PWM_STRETCH_VALUE7(0)
        , .PWM_STRETCH_VALUE8(0), .PWM_STRETCH_VALUE9(0), .SHADOW_REG_EN1(0)
        , .SHADOW_REG_EN10(0), .SHADOW_REG_EN11(0), .SHADOW_REG_EN12(0)
        , .SHADOW_REG_EN13(0), .SHADOW_REG_EN14(0), .SHADOW_REG_EN15(0)
        , .SHADOW_REG_EN16(0), .SHADOW_REG_EN2(0), .SHADOW_REG_EN3(0)
        , .SHADOW_REG_EN4(0), .SHADOW_REG_EN5(0), .SHADOW_REG_EN6(0), .SHADOW_REG_EN7(0)
        , .SHADOW_REG_EN8(0), .SHADOW_REG_EN9(0), .TACHINT_ACT_LEVEL(0)
        , .TACH_EDGE1(0), .TACH_EDGE10(0), .TACH_EDGE11(0), .TACH_EDGE12(0)
        , .TACH_EDGE13(0), .TACH_EDGE14(0), .TACH_EDGE15(0), .TACH_EDGE16(0)
        , .TACH_EDGE2(0), .TACH_EDGE3(0), .TACH_EDGE4(0), .TACH_EDGE5(0)
        , .TACH_EDGE6(0), .TACH_EDGE7(0), .TACH_EDGE8(0), .TACH_EDGE9(0)
        , .TACH_NUM(1) )  corepwm_0 (.PCLK(final_mss_0_FAB_CLK), 
        .PENABLE(CoreAPB3_0_APBmslave0_PENABLE), .PRESETN(
        final_mss_0_M2F_RESET_N), .PSEL(CoreAPB3_0_APBmslave0_PSELx), 
        .PREADY(CoreAPB3_0_APBmslave0_PREADY), .PSLVERR(
        CoreAPB3_0_APBmslave0_PSLVERR), .TACHINT(), .PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .PADDR({
        \CoreAPB3_0_APBmslave0_PADDR_[7] , 
        \CoreAPB3_0_APBmslave0_PADDR_[6] , 
        \CoreAPB3_0_APBmslave0_PADDR_[5] , 
        \CoreAPB3_0_APBmslave0_PADDR_[4] , 
        \CoreAPB3_0_APBmslave0_PADDR_[3] , 
        \CoreAPB3_0_APBmslave0_PADDR_[2] , 
        \CoreAPB3_0_APBmslave0_PADDR_[1] , 
        \CoreAPB3_0_APBmslave0_PADDR_[0] }), .PRDATA({
        \CoreAPB3_0_APBmslave0_PRDATA_[31] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PRDATA_[0] }), .PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA_[31] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[30] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[29] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[28] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[27] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[26] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[25] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[24] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[23] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[22] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[21] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[20] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[19] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[18] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[17] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[16] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[15] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[14] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[13] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[12] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[11] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[10] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[9] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[8] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] }), .TACHIN({TACHIN[1]}), 
        .PWM({PWM[8], PWM[7], PWM[6], PWM[5], PWM[4], PWM[3], PWM[2], 
        PWM[1]}));
    GND GND (.Y(GND_net));
    final_mss final_mss_0 (.MSS_RESET_N(MSS_RESET_N), .MSSPSEL(
        final_mss_0_MSS_MASTER_APB_PSELx), .MSSPENABLE(
        final_mss_0_MSS_MASTER_APB_PENABLE), .MSSPWRITE(
        final_mss_0_MSS_MASTER_APB_PWRITE), .MSSPREADY(
        final_mss_0_MSS_MASTER_APB_PREADY), .MSSPSLVERR(
        final_mss_0_MSS_MASTER_APB_PSLVERR), .M2F_RESET_N(
        final_mss_0_M2F_RESET_N), .UART_0_TXD(UART_0_TXD), .UART_0_RXD(
        UART_0_RXD), .FAB_CLK(final_mss_0_FAB_CLK), .ADCDirectInput_0(
        ADCDirectInput_0), .VAREF1(VAREF1), .UART_1_TXD(UART_1_TXD), 
        .UART_1_RXD(UART_1_RXD), .GPIO_15_OUT(GPIO_15_OUT), .MSSPADDR({
        \final_mss_0_MSS_MASTER_APB_PADDR_[19] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[18] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[17] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[16] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[15] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[14] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[13] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[12] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[11] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[10] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[9] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[8] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[7] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[6] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[5] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[4] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[3] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[2] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[1] , 
        \final_mss_0_MSS_MASTER_APB_PADDR_[0] }), .MSSPRDATA({
        \final_mss_0_MSS_MASTER_APB_PRDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PRDATA_[0] }), .MSSPWDATA({
        \final_mss_0_MSS_MASTER_APB_PWDATA_[31] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[30] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[29] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[28] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[27] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[26] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[25] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[24] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[23] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[22] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[21] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[20] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[19] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[18] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[17] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[16] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[15] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[14] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[13] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[12] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[11] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[10] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[9] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[8] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[7] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[6] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[5] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[4] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[3] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[2] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[1] , 
        \final_mss_0_MSS_MASTER_APB_PWDATA_[0] }));
    final_top_CoreUARTapb_0_CoreUARTapb #( .BAUD_VALUE(4800), .BAUD_VAL_FRCTN(0)
        , .BAUD_VAL_FRCTN_EN(0), .FAMILY(18), .FIXEDMODE(0), .PRG_BIT8(1)
        , .PRG_PARITY(0), .RX_FIFO(1), .RX_LEGACY_MODE(0), .TX_FIFO(1)
         )  CoreUARTapb_0 (.PCLK(final_mss_0_FAB_CLK), .PRESETN(
        final_mss_0_M2F_RESET_N), .PSEL(CoreAPB3_0_APBmslave2_PSELx), 
        .PENABLE(CoreAPB3_0_APBmslave0_PENABLE), .PWRITE(
        CoreAPB3_0_APBmslave0_PWRITE), .TXRDY(), .RXRDY(), .PARITY_ERR(
        ), .OVERFLOW(), .RX(RX), .TX(TX), .PREADY(
        CoreAPB3_0_APBmslave2_PREADY), .PSLVERR(
        CoreAPB3_0_APBmslave2_PSLVERR), .FRAMING_ERR(), .PADDR({
        \CoreAPB3_0_APBmslave1_PADDR_[4] , 
        \CoreAPB3_0_APBmslave1_PADDR_[3] , 
        \CoreAPB3_0_APBmslave1_PADDR_[2] , 
        \CoreAPB3_0_APBmslave1_PADDR_[1] , 
        \CoreAPB3_0_APBmslave1_PADDR_[0] }), .PWDATA({
        \CoreAPB3_0_APBmslave0_PWDATA_[7] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[6] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[5] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[4] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[3] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[2] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[1] , 
        \CoreAPB3_0_APBmslave0_PWDATA_[0] }), .PRDATA({
        \CoreAPB3_0_APBmslave2_PRDATA_[7] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[6] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[5] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[4] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[3] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[2] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[1] , 
        \CoreAPB3_0_APBmslave2_PRDATA_[0] }));
    
endmodule
